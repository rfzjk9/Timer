module alarm(rst,SW,sign,light,clk);
	input sign,rst,SW,clk;
	output reg[23:0] light;
	reg[4:0] i;
	always @(posedge clk) begin
	if(~rst) begin
		i = 0; end
	else
		if(SW) begin
			if(sign)	begin
				if(i<25) i = i+1;
				else i = 0;
				end
			else i = 0;
			end
		else i=0;
	end
	
	always @(i)
	case(i)
		0:light <= 24'b0000_0000_0000_0000_0000_0000;
		1:light <= 24'b1000_0000_0000_0000_0000_0000;
		2:light <= 24'b0100_0000_0000_0000_0000_0000;
		3:light <= 24'b0010_0000_0000_0000_0000_0000;
		4:light <= 24'b0001_0000_0000_0000_0000_0000;
		5:light <= 24'b0000_1000_0000_0000_0000_0000;
		6:light <= 24'b0000_0100_0000_0000_0000_0000;
		7:light <= 24'b0000_0010_0000_0000_0000_0000;
		8:light <= 24'b0000_0001_0000_0000_0000_0000;
		9:light <= 24'b0000_0000_1000_0000_0000_0000;
		10:light <= 24'b0000_0000_0100_0000_0000_0000;
		11:light <= 24'b0000_0000_0010_0000_0000_0000;
		12:light <= 24'b0000_0000_0001_0000_0000_0000;
		13:light <= 24'b0000_0000_0000_1000_0000_0000;
		14:light <= 24'b0000_0000_0000_0100_0000_0000;
		15:light <= 24'b0000_0000_0000_0010_0000_0000;
		16:light <= 24'b0000_0000_0000_0001_0000_0000;
		17:light <= 24'b0000_0000_0000_0000_1000_0000;
		18:light <= 24'b0000_0000_0000_0000_0100_0000;
		19:light <= 24'b0000_0000_0000_0000_0010_0000;
		20:light <= 24'b0000_0000_0000_0000_0001_0000;
		21:light <= 24'b0000_0000_0000_0000_0000_1000;
		22:light <= 24'b0000_0000_0000_0000_0000_0100;
		23:light <= 24'b0000_0000_0000_0000_0000_0010;
		24:light <= 24'b0000_0000_0000_0000_0000_0001;
		endcase
endmodule
